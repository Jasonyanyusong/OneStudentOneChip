//创建一个Verilog模块，实现与门的逻辑功能，如下图所示：
module top_module(
  input a, 
  input b,
  output out );
// 请用户在下方编辑代码
    assign out = a && b;
	
//用户编辑到此为止
endmodule
