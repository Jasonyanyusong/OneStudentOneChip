//编写 Verilog 代码，使电路输出信号0
module top_module(
  output out
);
  // Write your code here
    assign out = 1'b0;
endmodule