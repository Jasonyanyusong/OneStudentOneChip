module test_our_cpp;
    initial begin
        $display("Hello World");
        $finish;
    end
endmodule
