module mux_2to1 ();