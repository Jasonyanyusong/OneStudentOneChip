//创建一个名为top_module的Verilog模块，实现非门的功能
module top_module( input in, output out );
// 请用户在下方编辑代码
    assign out = !in;
  
//用户编辑到此为止
endmodule